ARCHITECTURE sim OF inverter IS
BEGIN

  out1 <= NOT in1;

END ARCHITECTURE sim;

